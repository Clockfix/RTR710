-- synopsis directives:
-- synthesis VHDL_INPUT_VERSION VHDL_2008

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

PACKAGE data_types IS
	TYPE aslv IS ARRAY(NATURAL RANGE <>) OF STD_LOGIC_VECTOR;
END PACKAGE;

PACKAGE BODY data_types IS
END PACKAGE BODY;